`define VERSION 0010